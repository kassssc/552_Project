module m(
	input branch_new,
	input memwrite_new,
	input memread_new,
	input clk,
	input rst, 
	input wen
);
