module CACHE (

);

endmodule